package IOCapAxi;

import IOCapAxi_Types :: *;
import IOCapAxi_Flits :: *;
import IOCapAxi_Exposers :: *;
import IOCapAxi_KeyManagers :: *;
import IOCapAxi_Windows :: *;

export IOCapAxi_Types :: *;
export IOCapAxi_Flits :: *;
export IOCapAxi_Exposers :: *;
export IOCapAxi_KeyManagers :: *;
export IOCapAxi_Windows :: *;

endpackage