(* synthesize *)
module mkSimpleIOCapKeyManager_Tb(Empty);
endmodule